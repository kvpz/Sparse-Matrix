100 2
200 2
300 2
1 2
799 2
